`define MODULE_NAME cic_filter
`define DECIMATOR
