`define MODULE_NAME integer_multiplier
`define SIGNED_A
`define SIGNED_B
`define DATA_B
`define LUT
`define NON_PIPELINE
