parameter DIN_WIDTH=32;
parameter M=2;
parameter N=4;
parameter R=177;
parameter DOUT_WIDTH=68;
parameter MODE=0;
