parameter WIDTH_B = 20;
parameter WIDTH_A = 12;
