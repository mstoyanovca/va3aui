`define DEFINE_FPGA_TYPE "GW1N"
`define DEFINE_WORKMODE 2
`define DEFINE_CH_NUM 1
`define DEFINE_PHASE_WIDTH 25
`define DEFINE_OUTPUT_WIDTH 20
`define DEFINE_PHASE_DITHER "NO"
`define DEFINE_TAYLOR_CORR "YES"
`define DEFINE_TRUNC_WIDTH 13
`define DEFINE_PINC_TYPE "Fixed"
`define DEFINE_POFF_TYPE "None"
`define PHASE_EN
`define PHASEIN_EN
`define SINE_OUT
`define COSSINE_OUT
`define DEFINE_DELAY 6
`define DEFINE_PINC0_INIT 25'h147AE1
`define DEFINE_POFF0_INIT 25'h0
`define DEFINE_PINC1_INIT 25'h0
`define DEFINE_POFF1_INIT 25'h0
`define DEFINE_PINC2_INIT 25'h0
`define DEFINE_POFF2_INIT 25'h0
`define DEFINE_PINC3_INIT 25'h0
`define DEFINE_POFF3_INIT 25'h0
`define DEFINE_PINC4_INIT 25'h0
`define DEFINE_POFF4_INIT 25'h0
`define DEFINE_PINC5_INIT 25'h0
`define DEFINE_POFF5_INIT 25'h0
`define DEFINE_PINC6_INIT 25'h0
`define DEFINE_POFF6_INIT 25'h0
`define DEFINE_PINC7_INIT 25'h0
`define DEFINE_POFF7_INIT 25'h0
`define DEFINE_PINC8_INIT 25'h0
`define DEFINE_POFF8_INIT 25'h0
`define DEFINE_PINC9_INIT 25'h0
`define DEFINE_POFF9_INIT 25'h0
`define DEFINE_PINCA_INIT 25'h0
`define DEFINE_POFFA_INIT 25'h0
`define DEFINE_PINCB_INIT 25'h0
`define DEFINE_POFFB_INIT 25'h0
`define DEFINE_PINCC_INIT 25'h0
`define DEFINE_POFFC_INIT 25'h0
`define DEFINE_PINCD_INIT 25'h0
`define DEFINE_POFFD_INIT 25'h0
`define DEFINE_PINCE_INIT 25'h0
`define DEFINE_POFFE_INIT 25'h0
`define DEFINE_PINCF_INIT 25'h0
`define DEFINE_POFFF_INIT 25'h0
`define DEFINE_FILENAME "cos_sin_lut.dat"
