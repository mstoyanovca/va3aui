`define module_name dds_top
