parameter DIN_WIDTH=32;
parameter M=1;
parameter N=3;
parameter R=89;
parameter DOUT_WIDTH=53;
parameter MODE=0;
