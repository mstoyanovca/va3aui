`define MODULE_NAME fir_hilbert
`define fir_type_hilbert
