parameter DIN_WIDTH = 16;
parameter COEFF_WIDTH = 18;
parameter DOUT_WIDTH = 16;
parameter NUM_CHN = 1;
parameter NUM_FACTOR = 2;
parameter TAPS_SIZE = 43;
parameter NUM_TDM = 1;
parameter COEFF_PATH = "./coeff.dat";
