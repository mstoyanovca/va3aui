`define module_name dds_ii
